`ifndef __AXI_TYPEDEF_SVH__
`define __AXI_TYPEDEF_SVH__

`define AXI_ADDR_WIDTH          32
`define AXI_ADDR_OFFSET         6
`define AXI_DATA_WIDTH          64
`define AXI_ID_WIDTH            4

`endif /* __AXI_TYPEDEF_SVH__ */
